module data_source_mux (
   input wire [31:0] wrdata_cpu,
	input wire [31:0] rddata_cpu,
	output reg [31:0] outdata
);

endmodule 