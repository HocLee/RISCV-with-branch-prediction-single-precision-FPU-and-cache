module mux_rddata(

);
endmodule 